use IEEE
